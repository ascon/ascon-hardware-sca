../../../LWC_rtl/LWC_SCA.vhd