../v2/Round.vhd