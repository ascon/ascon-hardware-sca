../v1/CryptoCore_SCA.vhd