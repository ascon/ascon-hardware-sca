../v3/LWC_config_32_3s.vhd