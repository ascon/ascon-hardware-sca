../v1/Round.vhd