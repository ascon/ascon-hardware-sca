../v1/LWC_config_32_2s.vhd